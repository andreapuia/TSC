/***********************************************************************
 * A SystemVerilog RTL model of an instruction regisgter
 *
 * An error can be injected into the design by invoking compilation with
 * the option:  +define+FORCE_LOAD_ERROR
 *
 **********************************************************************/

//functie -> timp de simulare 0
//task - > contine timp de simulare 

module instr_register
import instr_register_pkg::*;  // pachetul instr_register_pkg -> declaram semnalele in el
(input  logic          clk,
 input  logic          load_en,
 input  logic          reset_n,
 input  operand_t      operand_a,
 input  operand_t      operand_b,
 input  operand_t      operand_c,
 input  opcode_t       opcode,
 input  address_t      write_pointer,
 input  address_t      read_pointer,
 output  result_t       result,
 output instruction_t  instruction_word // DE AICI SE GENEREAZA SEMNALUL instruction_t CARE VA FI FOLOSIT IN INTERFATA
);
 // timeunit 1ns/1ns;

  instruction_t  iw_reg [0:31];  // an array of instruction_word structures // 2 la 32 operatii 
  
  //aici avem operatiile din instr_register_pkg

  // write to the register
  always@(posedge clk, negedge reset_n)   // write into register
    if (!reset_n) begin
      foreach (iw_reg[i]) //pentru fiecare valoare din array
        iw_reg[i] = '{opc:ZERO,default:0};  // reset to all zeros
    end
    else if (load_en) begin
      @(operand_a, operand_b, operand_c);
      case (opcode)
              //iw_reg[write_pointer] = '{opcode,operand_a,operand_b};
      ZERO  : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c, 'b0};
      PASSA : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c, operand_a};
      PASSB : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c,operand_b};
      ADD   : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c,$signed(operand_a + operand_b + operand_c)};
      SUB   : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c,$signed(operand_a - operand_b)};
      MULT  : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c,$signed(operand_a * operand_b)};
      DIV   : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c,$signed(operand_a / operand_b)};
      MOD   : iw_reg[write_pointer] = '{opcode, operand_a, operand_b, operand_c,$signed(operand_a % operand_b)};
    default : iw_reg[write_pointer] = '{opcode, operand_a, operand_b,  operand_c, 'x};
    endcase
    result = iw_reg[write_pointer].result;
  end
  
  // read from the register
  assign instruction_word = iw_reg[read_pointer];  // continuously read from register

// compile with +define+FORCE_LOAD_ERROR to inject a functional bug for verification to catch
`ifdef FORCE_LOAD_ERROR
initial begin
  force operand_b = operand_a; // cause wrong value to be loaded into operand_b
end
`endif

endmodule: instr_register
